module DataPath ( 
			input ir_on_adr, pc_on_adr, // address bus control
			input dbus_on_data, data_on_dbus, // data bus control
			input ld_ir, ld_ac, ld_pc, inc_pc, clr_pc, // ir and pc control
			input pass, add, // alu control
			input alu_on_dbus,
			input clk,
				
			output [5:0] adr_bus, // address bus out
			output [1:0] op_code, // first 2 bits of IR 
			inout [7:0] data_bus
);
				
	wire [7:0] dbus, ir_out, a_out, alu_out; // dbus - internal data bus
	wire [5:0] pc_out;
	
	IR ir (.data_in(dbus), 
			 .load(ld_ir), 
			 .clk(clk), 
			 .data_out(ir_out));
			 
	PC pc (.data_in(ir_out[5:0]), 
			 .load(ld_pc), .inc(inc_pc), 
			 .clr(clr_pc), 
			 .clk(clk), 
			 .data_out(pc_out));
			 
	AC ac (.data_in(dbus), 
			 .load(ld_ac),
			 .clk(clk),
			 .data_out(a_out)); 
 
 
	ALU alu (.a(a_out),
				.b({2'b00,ir_out[5:0]}),
				.pass(pass),
				.add(add),
				.alu_out(alu_out));
				
			

	assign adr_bus = ir_on_adr ? ir_out[5:0] : 6'bzz_zzzz; // ir to addr bus for jump instruction
	assign adr_bus = pc_on_adr ? pc_out : 6'bzz_zzzz; // pc to addr bus to fetch next instruction
	
	assign dbus = alu_on_dbus ? alu_out : 8'bzzzz_zzzz; // if alu result available, put it on internal data bus
	assign data_bus = dbus_on_data ? dbus : 8'bzzzz_zzzz; // internal to external data bus
	
	assign dbus = data_on_dbus ? data_bus : 8'bzzzz_zzzz; // if data available from external data bus, put it on internal
	
	assign op_code = ir_out[7:6]; // first 2 bits of IR
 
 
 endmodule